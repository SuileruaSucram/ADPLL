//Author: Jisu


//C stands for control signals
//F stands for frequencies

//todo: implement a register that convert 1 channal I2C bursts to 32bits

`timescale 1ps/1ps
module ADPLL(En, volt_0, volt_1, Reset,F_input,C_info,C_target, F_xtal,F_output1,F_output2);
	input En,Reset, volt_0, volt_1;		// enable, Reset
	input C_info;			//information whether the target is frequency(1) or multipler(0)
	input F_input;			//input frequency
	input [31:0]C_target;		//target frequency or multiplier which has one channel input with bursts of data (I2C)
	input F_xtal;			//Crystal oscillator : 50mhz
	output reg F_output1,F_output2; 

	wire [31:0] C_F2M1, C_F2M2;
	wire [31:0] C_N,C_1,C_2;
	wire [31:0] C_N1,C_N2;//controller output 
	
	wire [31:0]C_XR,C_RI;
	wire F_ring;			//frequency generated by the ring oscillator
	//module Ring (Clk, F_ring);
	Ring RingGenerate(F_input, volt_0, volt_1, F_ring);
	//module Freq_ratio(En,Reset,F_clk,F_ring,C_freq);
	Freq_ratioA Crystal_Input(En,Reset,F_xtal,F_ring,C_XR);

	Freq_ratioA Ring_Input(En,Reset,F_input,F_ring,C_RI);
	//assign C_RI = 32'd500000;
	
	//module Multiple_Calculator (En, Reset,Clk, Ratio_Crystal, Target_Freq, Multiplier);
	
	//Multiple_Calculator FreqToMulti(En, Reset,F_xtal, C_XI, C_target, C_F2M);
	
	//module Controller (En, Reset, C_N, C_Freq, C_N1, C_N2);
	Controller Process(En, Reset, C_target, C_RI, C_N1, C_N2);	
	//module TargetController (En, Reset, C_RX, C_N, C_N1,C_N2);
	TargetController Process2 (En, Reset, C_XR, C_target, C_F2M1, C_F2M2);

	//assign C_1 = (C_info)? C_N1:C_F2M1;
	//assign C_2 = (C_info)? C_N2:C_F2M2;
	
	//This below does not work as a mux, but we have identified that this is
	//Where the problem is. put Control signals directly into Divider to test
	//TargetController needs tuned.
	
	genvar i;
	generate 
	for (i = 0; i < 32; i++)
	begin : assign_C
			assign C_1[i] = (!C_info & C_N1[i]) | (C_info & C_F2M1[i]);
			assign C_2[i] = (!C_info & C_N2[i]) | (C_info & C_F2M2[i]);

	end
	endgenerate

	//module Divider(En,Reset,C_N,F_input,F_output);
	Divider first (En,Reset,C_1,F_ring,F_output1);
	
	Divider second(En,Reset,C_2,F_ring,F_output2);
	
	
	endmodule
	
	
	`timescale 1ps/1ps
module ADPLL_TB;

	reg En,Reset, volt_0, volt_1;		// enable, Reset
	reg C_info;			//information whether the target is frequency(1) or multipler(0)
	reg F_input;			//input frequency
	reg [31:0]C_target;		//target frequency or multiplier which has one channel input with bursts of data (I2C)
	reg F_xtal;			//Crystal oscillator : 50mhz
	wire F_output1,F_output2; 
	logic F_Exp1, F_Exp2;
	
//module ADPLL(En,Reset,F_input,C_info,C_target, F_xtal,F_output1,F_output2);
	ADPLL DUT (En, volt_0, volt_1, Reset,F_input,C_info,C_target, F_xtal,F_output1,F_output2);
always begin
	F_Exp1 =1'b0;
	#166666;
	F_Exp1 =1'b1;
	#166666;

end
always begin
	F_Exp2 = 1'b0;
	#250000;
	F_Exp2 = 1'b1;
	#250000;
end
always begin  	//crystal frequency is 50mhz
		F_xtal = 1'b0;  	
		#10000;  	
		F_xtal = 1'b1;  	
		#10000;  
	end 
always begin //input frequency is 1mhz
	F_input = 1;
	#500000;
	F_input = 0;
	#500000;
	end
initial begin
 
	En = 0;
	volt_0 = 0;
	volt_1 = 0;
	Reset = 1;
	C_info = 0; //Freq
	C_target = 32'b00000001000000000000000110000000;//2 and 3
	//         32'b000000000 0000000 000000000 0000000
	#1ns;
	Reset = 0;
	#1ns;
	En = 1;
	volt_0 = 1;
	volt_1 = 1;
	#0.3ms; // freq_ratio module aleast needs 100 cylcles of input frequency to get the output: 100*1/10^6 = 1* 10^-3
	$stop;

end

endmodule
	